/*	
*	Author:	Kayleigh Humphrey
*	Date: 	Oct. 10, 2023
*	Name:   	Next State Logic
*  Next State Logic equations obtained through K-maps from the State Transition Table.
*
*	Inputs:	
*	S[0], S[1], S[2] & S[3] - States
*	Y[0] & Y[1] - the encoded inputs, to be called in the top level
*	
*	Outputs:
*	D[0], D[1], D[2] & D[3] - Next State Logic Equations
*	
*/ 


module statelogic(
	input logic s[3:0],
	input logic y[1:0], 
	output logic d[3:0]
);

//assign d[0] = ((~s[1] & ~s[0] & ~y[1] &  y[0] & ~s[2] & ~s[3]) | (~s[1] & s[0] & ~y[1] & ~y[0] & ~s[2]& ~s[3]) | (~s[1] & s[0] & y[1] & ~s[2] & ~s[3])| (s[1] & s[0] & ~y[1] & y[0] & ~s[2] & ~s[3]) | (s[1] & ~s[0] & ~y[1] & ~y[0] & ~s[2] & ~s[3]) | (s[1] & ~s[0] & y[1] & ~s[2] & ~s[3]) | (~y[1] & y[0] & s[2] & ~s[3]) | (~s[1] & ~s[0] & y[0] & ~s[2] & s[3]));
//assign d[1] = ((~s[1] &  y[1] &  y[0] & ~s[2] & ~s[3]) | (~s[1] & s[0] & ~y[1] & y[0] & ~s[2] & ~s[3])| (s[1] & ~y[1] & ~y[0] & ~s[2] & ~s[3]) | (s[1] & ~s[0] & y[0] & ~s[2] & ~s[3]) | (s[1] & ~s[0] & y[1] & y[0] & ~s[2] & ~s[3]) | (y[1] & ~y[0] & s[2] & ~s[3]) | (~s[1] & ~s[0] & y[1] & ~s[2] & s[3]));
//assign d[2] = ((~s[3] & ~s[2] &  y[1] &  y[0]) | (~s[2] & ~s[3] & y[0] & s[1] & s[0]) | (~s[2] & ~s[3] & y[1] & s[1]) | (s[2] & ~s[3] & ~s[1] & ~s[0] & ~y[1]) | (s[2] & ~s[3] & ~s[1] & ~s[0] & y[1] & ~y[0]) | (s[2] & ~s[3] & y[1] & y[0] & s[0]) | (s[2] & ~s[3] & y[1] & y[0] & s[1]));
//assign d[3] = (( s[2] & ~s[3] &  y[1] &  y[0] & ~s[1] & ~s[0]));

assign d[0] = ((y[0] & ~y[1] & ~s[0] & ~s[1] & ~s[2] & ~s[3] ) | (~y[0] & ~y[1] & s[0] & ~s[2] & ~s[3]) | ( y[1] & s[0] & ~s[2] & ~s[3]) | (y[0] & ~y[1] & ~s[0] & s[1] & ~s[2] & ~s[3]) | (y[0] & ~y[1]  & ~s[1] & s[2] & ~s[3]) | (y[0] & ~y[1] & s[0] & s[1] & s[2] & ~s[3]) | ( y[1] & ~s[0] & s[1] & s[2] & ~s[3]) | ( y[1] & ~s[0] & ~s[1] & ~s[2] & s[3]));
assign d[1] = ((y[0] & ~y[1] & s[0] & ~s[1] & ~s[2] & ~s[3]) | (~y[0] & y[1] & ~s[1] & ~s[2] & ~s[3]) | (~y[0] & ~y[1] & s[1] & ~s[2] & ~s[3]) | (~y[1] & ~s[0] & s[1] & ~s[2] & ~s[3]) | (y[0] & ~s[0] & s[1] & ~s[2] & ~s[3]) | (y[0] & y[1] & s[1] & ~s[2] & ~s[3]) | (y[0] & ~y[1] & s[1] & s[2] & ~s[3]) | (y[0] & s[0] & s[1] & s[2] & ~s[3]) | (~y[0] & y[1] & ~s[1] & s[2] & ~s[3]) | (~y[0] & y[1] & ~s[0] & s[1] & s[2] & ~s[3]) | (y[0] & y[1] & ~s[0] & ~s[1] & ~s[2] & s[3]));
assign d[2] = ((y[0] & y[1] & ~s[2] & ~s[3] & ~s[1]) | (y[0] & s[0] & s[1] & ~s[2] & ~s[3]) | (y[1] & s[1] & ~s[2] & ~s[3]) | (~y[1] & ~s[0] & ~s[1] & s[2] & ~s[3]) | (~y[0] & ~s[0] & ~s[1] & s[2] & ~s[3]) |(y[0] & y[1] & s[0] & s[2] & ~s[3] ) | (y[1] & s[0] & s[1] & s[2] & ~s[3] ) | (y[0] & y[1] & s[1] & s[2] & ~s[3] ) | (y[0] & ~s[0] & ~s[1] & ~s[2] & s[3] ) | (y[1] & ~s[0] & ~s[1] & ~s[2] & s[3] ));
assign d[3] = ((y[0] & y[1] & ~s[0] & ~s[1] & s[2] & ~s[3]));

endmodule